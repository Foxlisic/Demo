/* verilator lint_off WIDTH */

module video
(
    input   wire        clock,
    output  reg [3:0]   r,
    output  reg [3:0]   g,
    output  reg [3:0]   b,
    output  wire        hs,
    output  wire        vs
);
// ---------------------------------------------------------------------
// Тайминги для горизонтальной и вертикальной развертки
parameter
//  Visible     Front       Sync        Back        Whole
    hzv =  640, hzf =   16, hzs =   96, hzb =   48, hzw =  800,
    vtv =  480, vtf =   10, vts =    2, vtb =   33, vtw =  525;
// ---------------------------------------------------------------------
assign hs = X < (hzb + hzv + hzf);
assign vs = Y < (vtb + vtv + vtf);
// ---------------------------------------------------------------------
wire        xmax = (X == hzw - 1);
wire        ymax = (Y == vtw - 1);
wire        show = X >= hzb && X < hzb+hzv && Y >= vtb && Y < vtb+vtv;
reg  [10:0] X    = 0;
reg  [10:0] Y    = 0;
wire [ 9:0] x    = X - hzb;
wire [ 9:0] y    = Y - vtb;
// ---------------------------------------------------------------------

// Окружность
wire    c1 = (x-320)*(x-320) + (y-240)*(y-240) < 100*100;               // Окружность
wire    c2 = (x-320)*(x-320) + (y-280)*(y-280) < 75*75 && (y < 280);    // Голова
wire    c3 = (x-280)*(x-280) + (y-255)*(y-255) < 8*8;                   // Левый и правый глаз
wire    c4 = (x-360)*(x-360) + (y-255)*(y-255) < 8*8;
wire    c5 = (x-250)*(x-250) + (y-200)*(y-200) < 6*6;   // Левое ухо
wire    c6 = (x-390)*(x-390) + (y-200)*(y-200) < 6*6;   // Правое ухо
wire    e1 = (x > y + 40)  && (x < y + 60)  && (x > 450 - y) && (y < 280);  // Левое ухо
wire    e2 = (x < 600 - y) && (x > 580 - y) && (x < y + 190) && (y < 280);  // Правое ухо
wire    g1 = (x[3:0] == 0 || y[3:0] == 0);                                  // Сетка
wire    s1 = ((x > 590 - y) && (x < y + 200) || (y > 280)) && (x + 35 > y); // Тень от лого

wire    xx = x[0] ^ y[0];

// Вывод видеосигнала
always @(posedge clock) begin

    // Кадровая развертка
    X <= xmax ?         0 : X + 1;
    Y <= xmax ? (ymax ? 0 : Y + 1) : Y;

    {r, g, b} <= 12'h000;

    // Вывод окна видеоадаптера
    if (X >= hzb && X < hzb+hzv && Y >= vtb && Y < vtb+vtv)
    begin
         {r, g, b} <=
            // Глаза
            c3 || c4 ? 12'h004 :
            // Андроид C2; C5:E1 левое; C6:E2 - правое ухо
            c2 || c5 || c6 || e1 || e2 ? 12'hFFF :
            // Фон кружок (сетка)
            c1 ? (s1 && xx ? 12'h000 : (g1 ? 12'h888 : 12'h047)) :
            // Фон общий
            12'hACC;
    end

end

endmodule
