/* verilator lint_off WIDTH */
module video
(
    input               clock,
    output  reg         r,
    output  reg         g,
    output  reg         b,
    output              hs,
    output              vs,
    input   [3:0]       key
);
// ---------------------------------------------------------------------
// Тайминги для горизонтальной и вертикальной развертки
parameter
//  Visible     Front       Sync        Back        Whole
    hzv =  640, hzf =   16, hzs =   96, hzb =   48, hzw =  800,
    vtv =  400, vtf =   12, vts =    2, vtb =   35, vtw =  449;
// ---------------------------------------------------------------------
assign hs = X < (hzb + hzv + hzf);
assign vs = Y < (vtb + vtv + vtf);
// ---------------------------------------------------------------------
reg  [ 9:0] X    = 0;
reg  [ 8:0] Y    = 0;
wire        xmax = (X == hzw - 1);
wire        ymax = (Y == vtw - 1);
wire        show = X >= hzb && X < hzb+hzv && Y >= vtb && Y < vtb+vtv;
// ---------------------------------------------------------------------
wire [ 5:0] G = {Y[2:0], X[2:0]};
wire [ 5:0] P =
    G == 8'h00 ? 0  : G == 8'h01 ? 32 : G == 8'h02 ?  8 : G == 8'h03 ? 40 :
    G == 8'h04 ?  2 : G == 8'h05 ? 34 : G == 8'h06 ? 10 : G == 8'h07 ? 42 :
    G == 8'h08 ? 48 : G == 8'h09 ? 16 : G == 8'h0A ? 56 : G == 8'h0B ? 24 :
    G == 8'h0C ? 50 : G == 8'h0D ? 18 : G == 8'h0E ? 58 : G == 8'h0F ? 26 :
    G == 8'h10 ? 12 : G == 8'h11 ? 44 : G == 8'h12 ? 4  : G == 8'h13 ? 36 :
    G == 8'h14 ? 14 : G == 8'h15 ? 46 : G == 8'h16 ? 6  : G == 8'h17 ? 38 :
    G == 8'h18 ? 60 : G == 8'h19 ? 28 : G == 8'h1A ? 52 : G == 8'h1B ? 20 :
    G == 8'h1C ? 62 : G == 8'h1D ? 30 : G == 8'h1E ? 54 : G == 8'h1F ? 22 :
    G == 8'h20 ? 3  : G == 8'h21 ? 35 : G == 8'h22 ? 11 : G == 8'h23 ? 43 :
    G == 8'h24 ? 1  : G == 8'h25 ? 33 : G == 8'h26 ? 9  : G == 8'h27 ? 41 :
    G == 8'h28 ? 51 : G == 8'h29 ? 19 : G == 8'h2A ? 59 : G == 8'h2B ? 27 :
    G == 8'h2C ? 49 : G == 8'h2D ? 17 : G == 8'h2E ? 57 : G == 8'h2F ? 25 :
    G == 8'h30 ? 15 : G == 8'h31 ? 47 : G == 8'h32 ? 7  : G == 8'h33 ? 39 :
    G == 8'h34 ? 13 : G == 8'h35 ? 45 : G == 8'h36 ? 5  : G == 8'h37 ? 37 :
    G == 8'h38 ? 63 : G == 8'h39 ? 31 : G == 8'h3A ? 55 : G == 8'h3B ? 23 :
    G == 8'h3C ? 61 : G == 8'h3D ? 29 : G == 8'h3E ? 53 : 21;

reg [16:0] rnd;
reg [7:0] K;

wire [7:0] x = X + K;

// Вывод видеосигнала
always @(posedge clock)
begin

    // Кадровая развертка
    X <= xmax ?         0 : X + 1;
    Y <= xmax ? (ymax ? 0 : Y + 1) : Y;
    K <= xmax && ymax ? K + 1 : K;

    {r, g, b} <= 3'b000;

    if (show) begin

        {r, g, b} <= 3'b011;

        rnd <= rnd ? (rnd >> 1) ^ {rnd[0], 2'b00, rnd[0], 13'b0} : 1'b1;

        // Окно
        if (X >= 150 && Y >= 100 && X < 600 && Y < 340) {r,g,b} <= 3'b000;
        if (X >= 151 && Y >= 101 && X < 599 && Y < 339) {r,g,b} <= 3'b111;
        if (X >= 152 && Y == 338 && X < 598) {r,g,b} <= 3'b000;
        if (X == 598 && Y >= 102 && Y < 339) {r,g,b} <= 3'b000;
        if (X >= 153 && X < 596 && Y >= 103 && Y <= 120) {r,g,b} <= ((X - 153) >> 3) < P ? 3'b001 : 3'b011;

        // Кнопка
        if (X >= 580 && Y >= 104 && X <= 594 && Y <= 119) {r,g,b} <= (X == 594 || Y == 119 || (X == 593 && Y[0]) || (Y == 118 && X[0]) || (X - 580 == Y - 104) || (13 - (X - 580) == Y - 104) ? 3'b000 : 3'b111);

        // DEMO
        if (X >= 153 && Y >= 122 && X < 421 && Y <= 336) {r,g,b} <= 3'b000;
        if (X >= 154 && Y >= 123 && X < 420 && Y <= 335) {r,g,b} <= rnd[2:0];

        // DEMO1
        if (X >= 423 && Y >= 122 && X < 597 && Y <= 336) {r,g,b} <= 3'b000;
        if (X >= 424 && Y >= 123 && X < 596 && Y <= 335) {r,g,b} <= (Y < 240 ? x[5:3] - Y[5:3] : x[5:3] ^ Y[5:3]);

    end

end

endmodule
